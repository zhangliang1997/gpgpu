import defines::*;

module fetch(
	input in,
	output logic out

);	


scalar_t  pcRegs[NUM_WRAPS_PER_CORE];
assign out = 1;

endmodule 

module fetch(

);	



endmodule 

package defines;

parameter NUM_WRAPS_PER_CORE 			= 4;
parameter NUM_CORES						= 2;

typedef  logic[31:0]  scalar_t;


endpackage : defines;

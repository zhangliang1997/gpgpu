package defines;

parameter NUM_WARPS_PER_SM  			= 4;
parameter NUM_SMS						= 2;

parameter RESET_PC                      = 0;

typedef  logic[31:0]  scalar_t;


endpackage

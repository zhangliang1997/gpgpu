import defines::*;

module ift_fetch_data(
	input logic clk,
	input logic reset,

	input  logic[L1I_TAG_WIDTH - 1 : 0]    tags[NUM_L1I_WAYS],
	input  logic							way_valid[NUM_L1I_WAYS]
);













endmodule 
